`ifndef PROGRAM_VENDING
`define PROGRAM_VENDING

parameter bit [31:0] INSTRUCTIONS_VENDING[0:45] = '{
  32'b00000011001000000000010000010011,
  32'b00000000010100000000010010010011,
  32'b00000000101000000000010100010011,
  32'b00000001100100000000010110010011,
  32'b00000000010000000010001100000011,
  32'b00000000000000000000001110010011,
  32'b01111111111100110111000100010011,
  32'b00000000001000100000001000110011,
  32'b00000100001000110001001001100011,
  32'b00000100000000101001001001100011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000010100000100101000001100011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000001010010011,
  32'b00000000011100000010010000100011,
  32'b00000000010000000010001100000011,
  32'b11111100010111111111000001101111,
  32'b10000000000000000000001110010011,
  32'b01000000100000100000001000110011,
  32'b00000000000100000000001010010011,
  32'b11111110100111111111000001101111,
  32'b00000000000100000000001010010011,
  32'b00000010101100100101000001100011,
  32'b00000010101000100101010001100011,
  32'b00000010100100100101100001100011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b11111100000000100000001011100011,
  32'b00000000000000000000000001110011,
  32'b00000000101100111110001110110011,
  32'b01000000101100100000001000110011,
  32'b00000001100000000000000001101111,
  32'b00000000101000111110001110110011,
  32'b01000000101000100000001000110011,
  32'b00000000110000000000000001101111,
  32'b00000000100100111110001110110011,
  32'b01000000100100100000001000110011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b11111000000000100000101011100011,
  32'b11111001010111111111000001101111
};

`endif