`ifndef CONSTANT_EXCEPTION
`define CONSTANT_EXCEPTION


`define INSTRUCTION_ADDRESS_MISALIGNED 0
`define INSTRUCTION_ACCESS_FAULT 1
`define ILLEGAL_INSTRUCTION 2
`define BREAKPOINT 3
`define LOAD_ADDRESS_MISALIGNED 4
`define LOAD_ACCESS_FAULT 5
`define STORE_ADDRESS_MISALIGNED 6
`define STORE_ACCESS_FAULT 7
`define ENVIRONMENT_CALL_FROM_UMODE 8
`define ENVIRONMENT_CALL_FROM_SMODE 9
`define ENVIRONMENT_CALL_FROM_MMODE 11
`define INSTRUCTION_PAGE_FAULT 12
`define LOAD_PAGE_FAULT 13
`define STORE_PAGE_FAULT 15
`define DOUBLE_TRAP 16
`define SOFTWARE_CHECK 18
`define HARDWARE_ERROR 19


`endif
