`ifndef PROGRAM_TEST
`define PROGRAM_TEST

parameter [31:0] INSTRUCTIONS_TEST[0:9] = {
  32'b00000000000000000000000100110111,
  32'b00000001001000010000000100010011,
  32'b00000000000000000000000110110111,
  32'b00000010010000011000000110010011,
  32'b00000000001100010000001000110011,
  32'b00000000001000000010000000100011,
  32'b00000000001100000010000000100011,
  32'b00000000010000000010000000100011,
  32'b00000000000100000000000001110011,
  32'b00000000000000000000000000010011
};

`endif