`ifndef PROGRAM_VENDING
`define PROGRAM_VENDING

parameter [31:0] INSTRUCTIONS_VENDING[0:35] = {
  32'b00000001111000000000010000010011,
  32'b00000000010100000000010010010011,
  32'b00000000101000000000010100010011,
  32'b00000000010000000010001100000011,
  32'b00000000111100110111000100010011,
  32'b00000000001000100000001000110011,
  32'b00000010100000100101110001100011,
  32'b00000000000000000000001110010011,
  32'b00000010001000110001110001100011,
  32'b00000010000000101001110001100011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000001010010011,
  32'b00000000011100000010010000100011,
  32'b00000000010000000010001100000011,
  32'b11111100010111111111000001101111,
  32'b00000001000000000000001110010011,
  32'b01000000100000100000001000110011,
  32'b00000000000100000000001010010011,
  32'b00000000101000100101110001100011,
  32'b00000010100100100101000001100011,
  32'b00000000000000000000000000010011,
  32'b00000000000000000000000000010011,
  32'b11111100000000100000101011100011,
  32'b00000000000000000000000001110011,
  32'b00000000101000111110001110110011,
  32'b01000000101000100000001000110011,
  32'b00000000110000000000000001101111,
  32'b00000000100100111110001110110011,
  32'b01000000100100100000001000110011,
  32'b11111010000000100000110011100011,
  32'b11111011100111111111000001101111
};

`endif